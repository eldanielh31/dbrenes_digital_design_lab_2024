module main(input  clock,
				input  reset,
				input logic direction,
				input logic moveH,
				input logic moveV,
				output [7:0] red,
				output [7:0] green,
				output [7:0] blue,
				output vgaclock,
				output hsync,
				output vsync,
				output n_blank);
				
				



endmodule 